module RAM #(
    parameter WIDTH = 16,
    parameter DEPTH = 15          
)(
    input  wire                 clk,
    input  wire                 load,
    input  wire [DEPTH-1:0] address,
    input  wire [WIDTH-1:0]     in,
    output wire [WIDTH-1:0]     out
);

    reg [WIDTH-1:0] mem [0:DEPTH-1];

    // écriture synchrone
    always @(posedge clk) begin
        if (load) begin
            mem[address] <= in;
        end
    end

    // lecture combinatoire
    assign out = mem[address];

endmodule
